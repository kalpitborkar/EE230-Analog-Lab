HW1 B4 RC Highpass filter

* Specifying the components
c1 1 2 0.1u
r1 2 0 10k

* Specifying the input voltage
vin 1 0 dc 0 ac 1 

.ac dec 10 1 1Meg
.control
run

* Plot Amplitude frequency response
plot vdb(2) xlog

.endc
.end