Half Wave precision rectifier

.include ua741.txt
.include Diode_1N914.txt

vin 1 0 sin(0 5 1k)
v1 3 0 -15
v2 4 0 15

x1 0 2 4 3 5 ua741
r1 1 2 10k
r2 2 6 10k
D1 2 5 1N914
D2 5 6 1N914

.tran 0.02ms 5ms
.control
run 

print v(1) v(5) v(6)

.endc 
.end

