Bridge Rectifier without capacitor

*Specifiying the input voltage
vin 1 0 sin(0 21.21 50)

* Including the 1N4007 diode model
.include 1N4007.spice.txt

* Specifying the diodes
D1 3 4 1N4007
D2 9 1 1N4007
D3 5 4 1N4007
D4 8 7 1N4007

* Specifying dummy voltages
vdummy1 1 3 0
vdummy2 8 9 0
vdummy3 0 5 0
vdummy4 7 0 0

* Specifying the load resistor
rL 4 8 500

* Specifying the capacitor
c1 4 8 1000u

.tran 0.01ms 300ms
.control
run

plot v(4) - v(8)
plot i(vdummy1) 
plot i(vdummy3)

.endc
.end


