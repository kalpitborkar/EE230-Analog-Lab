HW1 B1 RC Integrator Case 1

* Specifying the components
r1 1 2 10k
c1 2 0 0.1u

* Specifying the input voltage
*Case 1
vin 1 0 pulse(0 5 0 0 0 10ms 20ms) 

.tran 0.01ms 100ms
.control
run

plot v(1) v(2)

.endc
.end

