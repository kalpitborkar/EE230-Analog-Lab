Astable Multivibrator

.include ua741.txt

v1 5 0 15
v2 6 0 -15

r0 2 3 50k 
r1 1 0 30k
r2 3 1 35k
c1 2 0 0.01u

x1 1 2 5 6 3 ua741 

.tran 0.001ms 10ms
.control 
run 

print v(2) v(3)

.endc 
.end