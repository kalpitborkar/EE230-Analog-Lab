HW5 Q2 B NTC

* .include lm324.txt
.include ua741.txt
.include Thermistor.txt

vin 1 0 5
v1 7 0 15
v2 8 0 -15
r1 1 3 300
r2 1 2 300
r3 3 0 300 
r4 3 5 2k
r5 5 6 10k
r6 4 0 10k
r7 2 4 2k

x1 4 5 7 8 5 ua741
x2 2 0 temp_val thermistor Ro = 300 alpha = 3548
v_temp_val temp_val 0 20


* .dc temp_terminal 20 30 0.1
.dc v_temp_val 20 30 0.1
.control

run 
plot v(3)-v(2)

.endc 
.end 



