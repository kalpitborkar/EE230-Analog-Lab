Lab 5 Q2 A

.include ua741.txt

v1 3 0 15
v2 4 0 -15
v3 9 0 15
v4 10 0 -15
v5 14 0 15
v6 15 0 -15 
vref 6 0 0

vi1 17 7 0
vi2 17 12 0
vcm 17 0 2

r1 11 2 10k 
r2 2 5 10k 
r3 16 1 10k 
r4 1 6 10k
r5 13 16 10k
r6 8 11 10k 
r10 8 13 2.21k

x1 1 2 3 4 5 ua741 
x2 7 8 9 10 11 ua741 
x3 12 13 14 15 16 ua741 

.dc vcm -2 2 0.1
.control 
run 

plot v(5)/(v(7)-v(12))

.endc 
.end 
