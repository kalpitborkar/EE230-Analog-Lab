HW1 B2 RC Differentiator Case 1

* Specifying the components
c1 1 2 0.1u
r1 2 0 10k

* Specifying the input voltage
* Case 1
vin 1 0 pulse(0 5 0 0 0 10ms 20ms)

.tran 0.01ms 100ms
.control
run

plot v(1) v(2)

.endc
.end