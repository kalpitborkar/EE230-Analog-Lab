HW4 Q2

.include ua741.txt

vin 1 0 dc 0 ac 0.5
v1 4 0 15
v2 5 0 -15
r1 1 2 10k 
rx1 1 3 10k 
rx2 3 6 10k 
c1 2 0 47n

x1 2 3 4 5 6 ua741 

.ac dec 10 1 1Meg
.control 
run 

* Gain plot
plot 20*log10(abs(ac.v(6)/v(1))) xlog 
* Phase plot
plot {57.29*vp(6)} xlog

.endc 
.end
