HW5 Q2 A PTC

.include Thermistor.txt

* x1 1 0 temp_val thermistor Ro = 5K alpha = 3548  
x1 1 0 temp_val thermistor Ro = 300 alpha = -3548  

vin 1 0 5
v_temp_val temp_val 0 0

.dc v_temp_val 0 100 0.1
.control
run

plot -v(1)/i(vin) 

.endc 
.end 
