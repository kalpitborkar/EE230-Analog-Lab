Lab 5 Q1 B

.include lm324.txt

r1 1 4 1.4Meg 
r2 2 3 13.7k 
r3 2 0 280
c1 1 4 3.3p 
c2 2 0 1u 
cj 1 0 11p 

x1 2 1 3 0 4 lm324 

vcc 3 0 5
vref 2 0 0.1

i1 1 0 1.5u ac 1


.ac dec 10 1 100Meg
.control 
run 

plot vdb(4) xlog
plot 20*log10(abs(ac.v(4))) xlog 
* plot 20*log10(abs(ac.v(2))) xlog 

.endc 
.end 

