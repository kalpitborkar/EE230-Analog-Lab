Single-pole Active High-pass Filter

.include ua741.txt

vin 1 0 dc 0 ac 1
ra 2 0 4.7k
ca 1 2 0.1u
r1 3 6 9.1k
r2 3 0 1k

v1 4 0 12
v2 5 0 -12

x1 2 3 4 5 6 ua741

.ac dec 10 1 1Meg
.control
run

plot vdb(6) xlog
plot {57.29*vp(2)} xlog


.endc 
.end 

