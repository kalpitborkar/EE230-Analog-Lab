HW4 Q3 B 

.include ua741.txt

vin 1 0 pulse(-5v 5v 0 0 0 0.5ms 1ms)
v1 3 0 15
v2 4 0 -15
r1 1 2 18k 
r2 2 5 1.5Meg 
c1 2 5 47n 

x1 0 2 3 4 5 ua741

.tran 0.005ms 110ms 100ms
.control 
run 

plot v(1) v(5) 

.endc 
.end 



